module helloworld();

$display("HELLO WORLD");

endmodule

